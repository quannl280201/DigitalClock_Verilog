module mod_N_counter_tb;
	reg clk = 0;
	reg mode;
	reg up;
	reg down;
endmodule
